library ieee;
use ieee.std_logic_1164.all;

entity UNIT_NAME is
    --port (
    --  x : in std_logic;
    --  y : in std_logic;
    --);
end entity UNIT_NAME;

architecture UNIT_NAME_behavior of UNIT_NAME is
begin
end architecture UNIT_NAME_behavior;
